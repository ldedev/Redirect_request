module models

struct Status {
pub:
	msg  string
	code string = '200'
}
